package px_ss_csr_pkg;

parameter int PS_PX_SKIP_CR         = 0;
parameter int PS_PX_INTERVAL_CR     = 1;
parameter int PS_PX_ADD_INTERVAL_CR = 2;
parameter int PS_LN_SKIP_CR         = 3;
parameter int PS_LN_INTERVAL_CR     = 4;
parameter int PS_LN_ADD_INTERVAL_CR = 5;

parameter int TOTAL_CSR_CNT         = 6;

endpackage
