package blc_csr_pkg;

parameter int BLC_MODE_CR    = 0;
parameter int BLC_CAL_STB_CR = 1;
parameter int BLC_MAN_BL_CR  = 2;

parameter int BLC_CUR_BL_SR  = 3;

parameter int TOTAL_CSR_CNT  = 4;

endpackage
