package lut_ctrl_csr_pkg;

parameter LUT_ORIG_PX_CR = 0;
parameter LUT_MOD_PX_CR  = 1;
parameter LUT_WR_STB_CR  = 2;

parameter TOTAL_CSR_CNT  = 3;

endpackage
