package bilinear_demosaicing_3x3_csr_pkg;

parameter int DEMOSAICING_EN_CR      = 0;
parameter int DEMOSAICING_PATTERN_CR = 1;

parameter int TOTAL_CSR_CNT          = 2;

endpackage
