package white_balance_corrector_csr_pkg;

parameter int WB_MODE_CR     = 0;
parameter int WB_CAL_STB_CR  = 1;
parameter int WB_MAN_SEL_CR  = 2;
parameter int WB_MAN_COEF_CR = 3;
parameter int WB_MAN_LOCK_CR = 4;

parameter int WB_CUR_COEF_SR = 5;

parameter int TOTAL_CSR_CNT  = 6;

endpackage
