package conv_2d_csr_pkg;

parameter int WR_STB_CR     = 0;
parameter int COEF_NUM_CR   = 1;
parameter int COEF_VAL_CR   = 2;

parameter int TOTAL_CSR_CNT = 3;

endpackage
