package median_filter_csr_pkg;

parameter int MED_FILT_EN_CR = 0;

parameter int TOTAL_CSR_CNT  = 1;

endpackage
