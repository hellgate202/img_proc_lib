package color_corrector_csr_pkg;

parameter int CC_COEF_LOCK_CR = 0;
parameter int CC_COEF_SEL_CR  = 1;
parameter int CC_COEF_CR      = 2;

parameter int TOTAL_CSR_CNT   = 3;

endpackage
