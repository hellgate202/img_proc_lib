package lut_rom_pkg;

parameter logic [9 : 0] INIT_DATA [1023 : 0] = {
  10'h0,
  10'h2d,
  10'h3d,
  10'h4a,
  10'h54,
  10'h5d,
  10'h65,
  10'h6c,
  10'h73,
  10'h79,
  10'h7f,
  10'h85,
  10'h8a,
  10'h8f,
  10'h94,
  10'h98,
  10'h9d,
  10'ha1,
  10'ha6,
  10'haa,
  10'hae,
  10'hb2,
  10'hb5,
  10'hb9,
  10'hbd,
  10'hc0,
  10'hc3,
  10'hc7,
  10'hca,
  10'hcd,
  10'hd0,
  10'hd4,
  10'hd7,
  10'hda,
  10'hdd,
  10'he0,
  10'he2,
  10'he5,
  10'he8,
  10'heb,
  10'hed,
  10'hf0,
  10'hf3,
  10'hf5,
  10'hf8,
  10'hfa,
  10'hfd,
  10'hff,
  10'h102,
  10'h104,
  10'h107,
  10'h109,
  10'h10b,
  10'h10d,
  10'h110,
  10'h112,
  10'h114,
  10'h116,
  10'h119,
  10'h11b,
  10'h11d,
  10'h11f,
  10'h121,
  10'h123,
  10'h125,
  10'h127,
  10'h12a,
  10'h12c,
  10'h12e,
  10'h130,
  10'h132,
  10'h133,
  10'h135,
  10'h137,
  10'h139,
  10'h13b,
  10'h13d,
  10'h13f,
  10'h141,
  10'h143,
  10'h144,
  10'h146,
  10'h148,
  10'h14a,
  10'h14c,
  10'h14d,
  10'h14f,
  10'h151,
  10'h153,
  10'h154,
  10'h156,
  10'h158,
  10'h15a,
  10'h15b,
  10'h15d,
  10'h15f,
  10'h160,
  10'h162,
  10'h164,
  10'h165,
  10'h167,
  10'h168,
  10'h16a,
  10'h16c,
  10'h16d,
  10'h16f,
  10'h170,
  10'h172,
  10'h173,
  10'h175,
  10'h177,
  10'h178,
  10'h17a,
  10'h17b,
  10'h17d,
  10'h17e,
  10'h180,
  10'h181,
  10'h183,
  10'h184,
  10'h185,
  10'h187,
  10'h188,
  10'h18a,
  10'h18b,
  10'h18d,
  10'h18e,
  10'h190,
  10'h191,
  10'h192,
  10'h194,
  10'h195,
  10'h197,
  10'h198,
  10'h199,
  10'h19b,
  10'h19c,
  10'h19d,
  10'h19f,
  10'h1a0,
  10'h1a2,
  10'h1a3,
  10'h1a4,
  10'h1a6,
  10'h1a7,
  10'h1a8,
  10'h1a9,
  10'h1ab,
  10'h1ac,
  10'h1ad,
  10'h1af,
  10'h1b0,
  10'h1b1,
  10'h1b3,
  10'h1b4,
  10'h1b5,
  10'h1b6,
  10'h1b8,
  10'h1b9,
  10'h1ba,
  10'h1bb,
  10'h1bd,
  10'h1be,
  10'h1bf,
  10'h1c0,
  10'h1c2,
  10'h1c3,
  10'h1c4,
  10'h1c5,
  10'h1c6,
  10'h1c8,
  10'h1c9,
  10'h1ca,
  10'h1cb,
  10'h1cc,
  10'h1ce,
  10'h1cf,
  10'h1d0,
  10'h1d1,
  10'h1d2,
  10'h1d4,
  10'h1d5,
  10'h1d6,
  10'h1d7,
  10'h1d8,
  10'h1d9,
  10'h1db,
  10'h1dc,
  10'h1dd,
  10'h1de,
  10'h1df,
  10'h1e0,
  10'h1e1,
  10'h1e2,
  10'h1e4,
  10'h1e5,
  10'h1e6,
  10'h1e7,
  10'h1e8,
  10'h1e9,
  10'h1ea,
  10'h1eb,
  10'h1ec,
  10'h1ee,
  10'h1ef,
  10'h1f0,
  10'h1f1,
  10'h1f2,
  10'h1f3,
  10'h1f4,
  10'h1f5,
  10'h1f6,
  10'h1f7,
  10'h1f8,
  10'h1f9,
  10'h1fb,
  10'h1fc,
  10'h1fd,
  10'h1fe,
  10'h1ff,
  10'h200,
  10'h201,
  10'h202,
  10'h203,
  10'h204,
  10'h205,
  10'h206,
  10'h207,
  10'h208,
  10'h209,
  10'h20a,
  10'h20b,
  10'h20c,
  10'h20d,
  10'h20e,
  10'h20f,
  10'h210,
  10'h211,
  10'h212,
  10'h213,
  10'h214,
  10'h215,
  10'h216,
  10'h217,
  10'h218,
  10'h219,
  10'h21a,
  10'h21b,
  10'h21c,
  10'h21d,
  10'h21e,
  10'h21f,
  10'h220,
  10'h221,
  10'h222,
  10'h223,
  10'h224,
  10'h225,
  10'h226,
  10'h227,
  10'h228,
  10'h229,
  10'h22a,
  10'h22b,
  10'h22c,
  10'h22d,
  10'h22d,
  10'h22e,
  10'h22f,
  10'h230,
  10'h231,
  10'h232,
  10'h233,
  10'h234,
  10'h235,
  10'h236,
  10'h237,
  10'h238,
  10'h239,
  10'h23a,
  10'h23b,
  10'h23b,
  10'h23c,
  10'h23d,
  10'h23e,
  10'h23f,
  10'h240,
  10'h241,
  10'h242,
  10'h243,
  10'h244,
  10'h245,
  10'h245,
  10'h246,
  10'h247,
  10'h248,
  10'h249,
  10'h24a,
  10'h24b,
  10'h24c,
  10'h24d,
  10'h24d,
  10'h24e,
  10'h24f,
  10'h250,
  10'h251,
  10'h252,
  10'h253,
  10'h254,
  10'h254,
  10'h255,
  10'h256,
  10'h257,
  10'h258,
  10'h259,
  10'h25a,
  10'h25a,
  10'h25b,
  10'h25c,
  10'h25d,
  10'h25e,
  10'h25f,
  10'h260,
  10'h260,
  10'h261,
  10'h262,
  10'h263,
  10'h264,
  10'h265,
  10'h266,
  10'h266,
  10'h267,
  10'h268,
  10'h269,
  10'h26a,
  10'h26b,
  10'h26b,
  10'h26c,
  10'h26d,
  10'h26e,
  10'h26f,
  10'h26f,
  10'h270,
  10'h271,
  10'h272,
  10'h273,
  10'h274,
  10'h274,
  10'h275,
  10'h276,
  10'h277,
  10'h278,
  10'h278,
  10'h279,
  10'h27a,
  10'h27b,
  10'h27c,
  10'h27c,
  10'h27d,
  10'h27e,
  10'h27f,
  10'h280,
  10'h280,
  10'h281,
  10'h282,
  10'h283,
  10'h284,
  10'h284,
  10'h285,
  10'h286,
  10'h287,
  10'h288,
  10'h288,
  10'h289,
  10'h28a,
  10'h28b,
  10'h28c,
  10'h28c,
  10'h28d,
  10'h28e,
  10'h28f,
  10'h28f,
  10'h290,
  10'h291,
  10'h292,
  10'h293,
  10'h293,
  10'h294,
  10'h295,
  10'h296,
  10'h296,
  10'h297,
  10'h298,
  10'h299,
  10'h299,
  10'h29a,
  10'h29b,
  10'h29c,
  10'h29c,
  10'h29d,
  10'h29e,
  10'h29f,
  10'h29f,
  10'h2a0,
  10'h2a1,
  10'h2a2,
  10'h2a2,
  10'h2a3,
  10'h2a4,
  10'h2a5,
  10'h2a5,
  10'h2a6,
  10'h2a7,
  10'h2a8,
  10'h2a8,
  10'h2a9,
  10'h2aa,
  10'h2ab,
  10'h2ab,
  10'h2ac,
  10'h2ad,
  10'h2ae,
  10'h2ae,
  10'h2af,
  10'h2b0,
  10'h2b0,
  10'h2b1,
  10'h2b2,
  10'h2b3,
  10'h2b3,
  10'h2b4,
  10'h2b5,
  10'h2b6,
  10'h2b6,
  10'h2b7,
  10'h2b8,
  10'h2b8,
  10'h2b9,
  10'h2ba,
  10'h2bb,
  10'h2bb,
  10'h2bc,
  10'h2bd,
  10'h2bd,
  10'h2be,
  10'h2bf,
  10'h2c0,
  10'h2c0,
  10'h2c1,
  10'h2c2,
  10'h2c2,
  10'h2c3,
  10'h2c4,
  10'h2c5,
  10'h2c5,
  10'h2c6,
  10'h2c7,
  10'h2c7,
  10'h2c8,
  10'h2c9,
  10'h2c9,
  10'h2ca,
  10'h2cb,
  10'h2cc,
  10'h2cc,
  10'h2cd,
  10'h2ce,
  10'h2ce,
  10'h2cf,
  10'h2d0,
  10'h2d0,
  10'h2d1,
  10'h2d2,
  10'h2d2,
  10'h2d3,
  10'h2d4,
  10'h2d5,
  10'h2d5,
  10'h2d6,
  10'h2d7,
  10'h2d7,
  10'h2d8,
  10'h2d9,
  10'h2d9,
  10'h2da,
  10'h2db,
  10'h2db,
  10'h2dc,
  10'h2dd,
  10'h2dd,
  10'h2de,
  10'h2df,
  10'h2df,
  10'h2e0,
  10'h2e1,
  10'h2e1,
  10'h2e2,
  10'h2e3,
  10'h2e3,
  10'h2e4,
  10'h2e5,
  10'h2e5,
  10'h2e6,
  10'h2e7,
  10'h2e7,
  10'h2e8,
  10'h2e9,
  10'h2e9,
  10'h2ea,
  10'h2eb,
  10'h2eb,
  10'h2ec,
  10'h2ed,
  10'h2ed,
  10'h2ee,
  10'h2ef,
  10'h2ef,
  10'h2f0,
  10'h2f1,
  10'h2f1,
  10'h2f2,
  10'h2f3,
  10'h2f3,
  10'h2f4,
  10'h2f5,
  10'h2f5,
  10'h2f6,
  10'h2f7,
  10'h2f7,
  10'h2f8,
  10'h2f8,
  10'h2f9,
  10'h2fa,
  10'h2fa,
  10'h2fb,
  10'h2fc,
  10'h2fc,
  10'h2fd,
  10'h2fe,
  10'h2fe,
  10'h2ff,
  10'h300,
  10'h300,
  10'h301,
  10'h301,
  10'h302,
  10'h303,
  10'h303,
  10'h304,
  10'h305,
  10'h305,
  10'h306,
  10'h307,
  10'h307,
  10'h308,
  10'h308,
  10'h309,
  10'h30a,
  10'h30a,
  10'h30b,
  10'h30c,
  10'h30c,
  10'h30d,
  10'h30d,
  10'h30e,
  10'h30f,
  10'h30f,
  10'h310,
  10'h311,
  10'h311,
  10'h312,
  10'h312,
  10'h313,
  10'h314,
  10'h314,
  10'h315,
  10'h315,
  10'h316,
  10'h317,
  10'h317,
  10'h318,
  10'h319,
  10'h319,
  10'h31a,
  10'h31a,
  10'h31b,
  10'h31c,
  10'h31c,
  10'h31d,
  10'h31d,
  10'h31e,
  10'h31f,
  10'h31f,
  10'h320,
  10'h321,
  10'h321,
  10'h322,
  10'h322,
  10'h323,
  10'h324,
  10'h324,
  10'h325,
  10'h325,
  10'h326,
  10'h327,
  10'h327,
  10'h328,
  10'h328,
  10'h329,
  10'h32a,
  10'h32a,
  10'h32b,
  10'h32b,
  10'h32c,
  10'h32d,
  10'h32d,
  10'h32e,
  10'h32e,
  10'h32f,
  10'h330,
  10'h330,
  10'h331,
  10'h331,
  10'h332,
  10'h332,
  10'h333,
  10'h334,
  10'h334,
  10'h335,
  10'h335,
  10'h336,
  10'h337,
  10'h337,
  10'h338,
  10'h338,
  10'h339,
  10'h33a,
  10'h33a,
  10'h33b,
  10'h33b,
  10'h33c,
  10'h33c,
  10'h33d,
  10'h33e,
  10'h33e,
  10'h33f,
  10'h33f,
  10'h340,
  10'h340,
  10'h341,
  10'h342,
  10'h342,
  10'h343,
  10'h343,
  10'h344,
  10'h345,
  10'h345,
  10'h346,
  10'h346,
  10'h347,
  10'h347,
  10'h348,
  10'h349,
  10'h349,
  10'h34a,
  10'h34a,
  10'h34b,
  10'h34b,
  10'h34c,
  10'h34d,
  10'h34d,
  10'h34e,
  10'h34e,
  10'h34f,
  10'h34f,
  10'h350,
  10'h350,
  10'h351,
  10'h352,
  10'h352,
  10'h353,
  10'h353,
  10'h354,
  10'h354,
  10'h355,
  10'h356,
  10'h356,
  10'h357,
  10'h357,
  10'h358,
  10'h358,
  10'h359,
  10'h359,
  10'h35a,
  10'h35b,
  10'h35b,
  10'h35c,
  10'h35c,
  10'h35d,
  10'h35d,
  10'h35e,
  10'h35e,
  10'h35f,
  10'h360,
  10'h360,
  10'h361,
  10'h361,
  10'h362,
  10'h362,
  10'h363,
  10'h363,
  10'h364,
  10'h365,
  10'h365,
  10'h366,
  10'h366,
  10'h367,
  10'h367,
  10'h368,
  10'h368,
  10'h369,
  10'h369,
  10'h36a,
  10'h36b,
  10'h36b,
  10'h36c,
  10'h36c,
  10'h36d,
  10'h36d,
  10'h36e,
  10'h36e,
  10'h36f,
  10'h36f,
  10'h370,
  10'h371,
  10'h371,
  10'h372,
  10'h372,
  10'h373,
  10'h373,
  10'h374,
  10'h374,
  10'h375,
  10'h375,
  10'h376,
  10'h376,
  10'h377,
  10'h378,
  10'h378,
  10'h379,
  10'h379,
  10'h37a,
  10'h37a,
  10'h37b,
  10'h37b,
  10'h37c,
  10'h37c,
  10'h37d,
  10'h37d,
  10'h37e,
  10'h37e,
  10'h37f,
  10'h380,
  10'h380,
  10'h381,
  10'h381,
  10'h382,
  10'h382,
  10'h383,
  10'h383,
  10'h384,
  10'h384,
  10'h385,
  10'h385,
  10'h386,
  10'h386,
  10'h387,
  10'h387,
  10'h388,
  10'h388,
  10'h389,
  10'h389,
  10'h38a,
  10'h38b,
  10'h38b,
  10'h38c,
  10'h38c,
  10'h38d,
  10'h38d,
  10'h38e,
  10'h38e,
  10'h38f,
  10'h38f,
  10'h390,
  10'h390,
  10'h391,
  10'h391,
  10'h392,
  10'h392,
  10'h393,
  10'h393,
  10'h394,
  10'h394,
  10'h395,
  10'h395,
  10'h396,
  10'h396,
  10'h397,
  10'h397,
  10'h398,
  10'h398,
  10'h399,
  10'h39a,
  10'h39a,
  10'h39b,
  10'h39b,
  10'h39c,
  10'h39c,
  10'h39d,
  10'h39d,
  10'h39e,
  10'h39e,
  10'h39f,
  10'h39f,
  10'h3a0,
  10'h3a0,
  10'h3a1,
  10'h3a1,
  10'h3a2,
  10'h3a2,
  10'h3a3,
  10'h3a3,
  10'h3a4,
  10'h3a4,
  10'h3a5,
  10'h3a5,
  10'h3a6,
  10'h3a6,
  10'h3a7,
  10'h3a7,
  10'h3a8,
  10'h3a8,
  10'h3a9,
  10'h3a9,
  10'h3aa,
  10'h3aa,
  10'h3ab,
  10'h3ab,
  10'h3ac,
  10'h3ac,
  10'h3ad,
  10'h3ad,
  10'h3ae,
  10'h3ae,
  10'h3af,
  10'h3af,
  10'h3b0,
  10'h3b0,
  10'h3b1,
  10'h3b1,
  10'h3b2,
  10'h3b2,
  10'h3b3,
  10'h3b3,
  10'h3b4,
  10'h3b4,
  10'h3b5,
  10'h3b5,
  10'h3b6,
  10'h3b6,
  10'h3b7,
  10'h3b7,
  10'h3b8,
  10'h3b8,
  10'h3b9,
  10'h3b9,
  10'h3ba,
  10'h3ba,
  10'h3bb,
  10'h3bb,
  10'h3bb,
  10'h3bc,
  10'h3bc,
  10'h3bd,
  10'h3bd,
  10'h3be,
  10'h3be,
  10'h3bf,
  10'h3bf,
  10'h3c0,
  10'h3c0,
  10'h3c1,
  10'h3c1,
  10'h3c2,
  10'h3c2,
  10'h3c3,
  10'h3c3,
  10'h3c4,
  10'h3c4,
  10'h3c5,
  10'h3c5,
  10'h3c6,
  10'h3c6,
  10'h3c7,
  10'h3c7,
  10'h3c8,
  10'h3c8,
  10'h3c9,
  10'h3c9,
  10'h3ca,
  10'h3ca,
  10'h3ca,
  10'h3cb,
  10'h3cb,
  10'h3cc,
  10'h3cc,
  10'h3cd,
  10'h3cd,
  10'h3ce,
  10'h3ce,
  10'h3cf,
  10'h3cf,
  10'h3d0,
  10'h3d0,
  10'h3d1,
  10'h3d1,
  10'h3d2,
  10'h3d2,
  10'h3d3,
  10'h3d3,
  10'h3d4,
  10'h3d4,
  10'h3d4,
  10'h3d5,
  10'h3d5,
  10'h3d6,
  10'h3d6,
  10'h3d7,
  10'h3d7,
  10'h3d8,
  10'h3d8,
  10'h3d9,
  10'h3d9,
  10'h3da,
  10'h3da,
  10'h3db,
  10'h3db,
  10'h3dc,
  10'h3dc,
  10'h3dd,
  10'h3dd,
  10'h3dd,
  10'h3de,
  10'h3de,
  10'h3df,
  10'h3df,
  10'h3e0,
  10'h3e0,
  10'h3e1,
  10'h3e1,
  10'h3e2,
  10'h3e2,
  10'h3e3,
  10'h3e3,
  10'h3e4,
  10'h3e4,
  10'h3e4,
  10'h3e5,
  10'h3e5,
  10'h3e6,
  10'h3e6,
  10'h3e7,
  10'h3e7,
  10'h3e8,
  10'h3e8,
  10'h3e9,
  10'h3e9,
  10'h3ea,
  10'h3ea,
  10'h3ea,
  10'h3eb,
  10'h3eb,
  10'h3ec,
  10'h3ec,
  10'h3ed,
  10'h3ed,
  10'h3ee,
  10'h3ee,
  10'h3ef,
  10'h3ef,
  10'h3f0,
  10'h3f0,
  10'h3f0,
  10'h3f1,
  10'h3f1,
  10'h3f2,
  10'h3f2,
  10'h3f3,
  10'h3f3,
  10'h3f4,
  10'h3f4,
  10'h3f5,
  10'h3f5,
  10'h3f5,
  10'h3f6,
  10'h3f6,
  10'h3f7,
  10'h3f7,
  10'h3f8,
  10'h3f8,
  10'h3f9,
  10'h3f9,
  10'h3fa,
  10'h3fa,
  10'h3fa,
  10'h3fb,
  10'h3fb,
  10'h3fc,
  10'h3fc,
  10'h3fd,
  10'h3fd,
  10'h3fe,
  10'h3fe,
  10'h3ff };

endpackage
